localparam position_01 = B1_51;
localparam position_02 = B1_16;
localparam position_03 = B1_35;
localparam position_04 = B1_08;
localparam position_05 = B1_34;
localparam position_06 = B1_36;
localparam position_07 = B1_12;
localparam position_08 = B1_44;
localparam position_09 = B1_31;
localparam position_10 = B1_03;
localparam position_11 = B1_32;
localparam position_12 = B1_01;
localparam position_13 = B1_49;
localparam position_14 = B1_07;
localparam position_15 = B1_20;
localparam position_16 = B1_42;
localparam position_17 = B1_47;
localparam position_18 = B1_26;
localparam position_19 = B1_39;
localparam position_20 = B1_46;
localparam position_21 = B1_02;
localparam position_22 = B1_13;
localparam position_23 = B1_24;
localparam position_24 = B1_40;
localparam position_25 = B1_11;
localparam position_26 = B1_33;
localparam position_27 = B1_38;
localparam position_28 = B1_23;
localparam position_29 = B1_10;
localparam position_30 = B1_45;
localparam position_31 = B1_04;
localparam position_32 = B1_29;
localparam position_33 = B1_27;
localparam position_34 = B1_18;
localparam position_35 = B1_37;
localparam position_36 = B1_28;
localparam position_37 = B1_09;
localparam position_38 = B1_21;
localparam position_39 = B1_52;
localparam position_40 = B1_30;
localparam position_41 = B1_05;
localparam position_42 = B1_22;
localparam position_43 = B1_43;
localparam position_44 = B1_48;
localparam position_45 = B1_14;
localparam position_46 = B1_50;
localparam position_47 = B1_41;
localparam position_48 = B1_25;
localparam position_49 = B1_17;
localparam position_50 = B1_19;
localparam position_51 = B1_15;
localparam position_52 = B1_06;